 /*                                                                      
 Copyright 2025 Haoyu Tang, haoyu.tang@hotmail.com
                                                                         
 Licensed under the Apache License, Version 2.0 (the "License");         
 you may not use this file except in compliance with the License.        
 You may obtain a copy of the License at                                 
                                                                         
     http://www.apache.org/licenses/LICENSE-2.0                          
                                                                         
 Unless required by applicable law or agreed to in writing, software    
 distributed under the License is distributed on an "AS IS" BASIS,       
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and     
 limitations under the License.                                          
 */

 module exu_alu_agu #(
    parameter A =1
 ) (
    input i_mem_wreq,
    input i_mem_rreq,
    input [31:0] i_alu_res,
    output o_mem_wen,
    output [31:0] o_mem_addr,
    output [31:0] o_mem_wdata,
    output o_mem_ren
 );

   assign o_mem_ren = i_mem_rreq;
   assign o_mem_wen = i_mem_wreq;
   assign o_mem_addr = i_alu_res;
    
 endmodule